    // *************************************************************
    // ASCII/Unicode Character ROM
    // *************************************************************

    module ascii_rom_th(
        input clk,
        input wire [10:0] addr,
        output reg [7:0] data
    );

    (* rom_style = "block" *) // Infer BRAM

    reg [10:0] addr_reg;

    always @(posedge clk)
        addr_reg <= addr;

    always @*
        case(addr_reg)
    
    // code x61 (ฟ)
        11'h610: data = 8'b00000001;	//        *
        11'h611: data = 8'b00000001;	//        *
        11'h612: data = 8'b00000001;	//        *
        11'h613: data = 8'b01101101;	//  ** ** *
        11'h614: data = 8'b00101101;	//   * ** *
        11'h615: data = 8'b01101101;	//  ** ** *
        11'h616: data = 8'b00110011;	//   **  **
        11'h617: data = 8'b00110011;	//   **  **
        11'h618: data = 8'b00110011;	//   **  **
        11'h619: data = 8'b00100001;	//   *    *
        11'h61a: data = 8'b00000000;	//         
        11'h61b: data = 8'b00000000;	//         
        11'h61c: data = 8'b00000000;	//         
        11'h61d: data = 8'b00000000;	//         
        11'h61e: data = 8'b00000000;	//         
        11'h61f: data = 8'b00000000;	//         

    // code x62 (ิ)
        11'he340: data = 8'b00000000;
        11'he341: data = 8'b00000000;
        11'he342: data = 8'b00000000;
        11'he343: data = 8'b00000000;
        11'he344: data = 8'b00111100;
        11'he345: data = 8'b01000010;
        11'he346: data = 8'b01111110;
        11'he347: data = 8'b00000000;
        11'he348: data = 8'b00000000;
        11'he349: data = 8'b00000000;
        11'he34a: data = 8'b00000000;
        11'he34b: data = 8'b00000000;
        11'he34c: data = 8'b00000000;
        11'he34d: data = 8'b00000000;
        11'he34e: data = 8'b00000000;
        11'he34f: data = 8'b00000000;

    // code x63 (แ)
        11'h630: data = 8'b00000000;	//         
        11'h631: data = 8'b00000000;	//         
        11'h632: data = 8'b00000000;	//         
        11'h633: data = 8'b01001000;	//  *  *   
        11'h634: data = 8'b01001000;	//  *  *   
        11'h635: data = 8'b01001000;	//  *  *   
        11'h636: data = 8'b01001000;	//  *  *   
        11'h637: data = 8'b01101100;	//  ** **  
        11'h638: data = 8'b01111110;	//  ****** 
        11'h639: data = 8'b01101100;	//  ** **  
        11'h63a: data = 8'b00000000;	//         
        11'h63b: data = 8'b00000000;	//         
        11'h63c: data = 8'b00000000;	//         
        11'h63d: data = 8'b00000000;	//         
        11'h63e: data = 8'b00000000;	//         
        11'h63f: data = 8'b00000000;	//         

    // code x64 (ก)
        11'h640: data = 8'b00000000;	//         
        11'h641: data = 8'b00000000;	//         
        11'h642: data = 8'b00000000;	//         
        11'h643: data = 8'b00111000;	//   ***   
        11'h644: data = 8'b01000100;	//  *   *  
        11'h645: data = 8'b01100100;	//  **  *  
        11'h646: data = 8'b01000100;	//  *   *  
        11'h647: data = 8'b01000100;	//  *   *  
        11'h648: data = 8'b01000100;	//  *   *  
        11'h649: data = 8'b01000100;	//  *   *  
        11'h64a: data = 8'b00000000;	//         
        11'h64b: data = 8'b00000000;	//         
        11'h64c: data = 8'b00000000;	//         
        11'h64d: data = 8'b00000000;	//         
        11'h64e: data = 8'b00000000;	//         
        11'h64f: data = 8'b00000000;	//         

    // code x65 (ำ)
        11'h650: data = 8'b00000000;	//         
        11'h651: data = 8'b00000000;	//         
        11'h652: data = 8'b00000000;	//         
        11'h653: data = 8'b01110000;	//  ***    
        11'h654: data = 8'b01001000;	//  *  *   
        11'h655: data = 8'b00001000;	//     *   
        11'h656: data = 8'b00001000;	//     *   
        11'h657: data = 8'b00001000;	//     *   
        11'h658: data = 8'b00001000;	//     *   
        11'h659: data = 8'b00001000;	//     *   
        11'h65a: data = 8'b00000000;	//         
        11'h65b: data = 8'b00000000;	//         
        11'h65c: data = 8'b00000000;	//         
        11'h65d: data = 8'b00000000;	//         
        11'h65e: data = 8'b00000000;	//         
        11'h65f: data = 8'b00000000;	//         

    // code x66 (ด)
        11'h660: data = 8'b00000000;	//         
        11'h661: data = 8'b00000000;	//         
        11'h662: data = 8'b00000000;	//         
        11'h663: data = 8'b01110000;	//  ***    
        11'h664: data = 8'b10001000;	// *   *   
        11'h665: data = 8'b10101000;	// * * *   
        11'h666: data = 8'b10101000;	// * * *   
        11'h667: data = 8'b10101000;	// * * *   
        11'h668: data = 8'b11001000;	// **  *   
        11'h669: data = 8'b11001000;	// **  *   
        11'h66a: data = 8'b00000000;	//         
        11'h66b: data = 8'b00000000;	//         
        11'h66c: data = 8'b00000000;	//         
        11'h66d: data = 8'b00000000;	//         
        11'h66e: data = 8'b00000000;	//         
        11'h66f: data = 8'b00000000;	//         

    // code x67 (เ)
        11'h670: data = 8'b00000000;	//         
        11'h671: data = 8'b00000000;	//         
        11'h672: data = 8'b00000000;	//         
        11'h673: data = 8'b01000000;	//  *      
        11'h674: data = 8'b01000000;	//  *      
        11'h675: data = 8'b01000000;	//  *      
        11'h676: data = 8'b01000000;	//  *      
        11'h677: data = 8'b01100000;	//  **     
        11'h678: data = 8'b01110000;	//  ***    
        11'h679: data = 8'b01100000;	//  **     
        11'h67a: data = 8'b00000000;	//         
        11'h67b: data = 8'b00000000;	//         
        11'h67c: data = 8'b00000000;	//         
        11'h67d: data = 8'b00000000;	//         
        11'h67e: data = 8'b00000000;	//         
        11'h67f: data = 8'b00000000;	//         

    // code x68 (้)
        11'h680: data = 8'b00000000;	//         
        11'h681: data = 8'b00000000;	//         
        11'h682: data = 8'b00000000;	//         
        11'h683: data = 8'b00000000;	//         
        11'h684: data = 8'b00000000;	//         
        11'h685: data = 8'b00000000;	//         
        11'h686: data = 8'b00000000;	//         
        11'h687: data = 8'b00000000;	//         
        11'h688: data = 8'b00000000;	//         
        11'h689: data = 8'b00000000;	//         
        11'h68a: data = 8'b00000000;	//         
        11'h68b: data = 8'b00000000;	//         
        11'h68c: data = 8'b00000000;	//         
        11'h68d: data = 8'b00000000;	//         
        11'h68e: data = 8'b00000000;	//         
        11'h68f: data = 8'b00000000;	//         

    // code x69 (ร)
        11'h690: data = 8'b00000000;	//         
        11'h691: data = 8'b00000000;	//         
        11'h692: data = 8'b00000000;	//         
        11'h693: data = 8'b11110000;	// ****    
        11'h694: data = 8'b11100000;	// ***     
        11'h695: data = 8'b00010000;	//    *    
        11'h696: data = 8'b00010000;	//    *    
        11'h697: data = 8'b00110000;	//   **    
        11'h698: data = 8'b00110000;	//   **    
        11'h699: data = 8'b00110000;	//   **    
        11'h69a: data = 8'b00000000;	//         
        11'h69b: data = 8'b00000000;	//         
        11'h69c: data = 8'b00000000;	//         
        11'h69d: data = 8'b00000000;	//         
        11'h69e: data = 8'b00000000;	//         
        11'h69f: data = 8'b00000000;	//         

    // code x6a (่)
        11'h6a0: data = 8'b11111111;	// ********
        11'h6a1: data = 8'b11111111;	// ********
        11'h6a2: data = 8'b11111111;	// ********
        11'h6a3: data = 8'b11111111;	// ********
        11'h6a4: data = 8'b11111111;	// ********
        11'h6a5: data = 8'b11111111;	// ********
        11'h6a6: data = 8'b11111111;	// ********
        11'h6a7: data = 8'b11111111;	// ********
        11'h6a8: data = 8'b11111111;	// ********
        11'h6a9: data = 8'b11111111;	// ********
        11'h6aa: data = 8'b11111111;	// ********
        11'h6ab: data = 8'b11111111;	// ********
        11'h6ac: data = 8'b11111111;	// ********
        11'h6ad: data = 8'b11111111;	// ********
        11'h6ae: data = 8'b11111111;	// ********
        11'h6af: data = 8'b11111111;	// ********

    // code x6b (า)
        11'h6b0: data = 8'b00000000;	//         
        11'h6b1: data = 8'b00000000;	//         
        11'h6b2: data = 8'b00000000;	//         
        11'h6b3: data = 8'b01110000;	//  ***    
        11'h6b4: data = 8'b01001000;	//  *  *   
        11'h6b5: data = 8'b00001000;	//     *   
        11'h6b6: data = 8'b00001000;	//     *   
        11'h6b7: data = 8'b00001000;	//     *   
        11'h6b8: data = 8'b00001000;	//     *   
        11'h6b9: data = 8'b00001000;	//     *   
        11'h6ba: data = 8'b00000000;	//         
        11'h6bb: data = 8'b00000000;	//         
        11'h6bc: data = 8'b00000000;	//         
        11'h6bd: data = 8'b00000000;	//         
        11'h6be: data = 8'b00000000;	//         
        11'h6bf: data = 8'b00000000;	//         

    // code x6c (ส)
        11'h6c0: data = 8'b00000000;	//         
        11'h6c1: data = 8'b00000000;	//         
        11'h6c2: data = 8'b00000100;	//      *  
        11'h6c3: data = 8'b00111100;	//   ****  
        11'h6c4: data = 8'b01001100;	//  *  **  
        11'h6c5: data = 8'b00110100;	//   ** *  
        11'h6c6: data = 8'b01101100;	//  ** **  
        11'h6c7: data = 8'b01000100;	//  *   *  
        11'h6c8: data = 8'b01100100;	//  **  *  
        11'h6c9: data = 8'b01100100;	//  **  *  
        11'h6ca: data = 8'b00000000;	//         
        11'h6cb: data = 8'b00000000;	//         
        11'h6cc: data = 8'b00000000;	//         
        11'h6cd: data = 8'b00000000;	//         
        11'h6ce: data = 8'b00000000;	//         
        11'h6cf: data = 8'b00000000;	//         

    // code x6d (ท)
        11'h6d0: data = 8'b00000000;	//         
        11'h6d1: data = 8'b00000000;	//         
        11'h6d2: data = 8'b00000000;	//         
        11'h6d3: data = 8'b01100110;	//  **  ** 
        11'h6d4: data = 8'b00101010;	//   * * * 
        11'h6d5: data = 8'b01101010;	//  ** * * 
        11'h6d6: data = 8'b00110010;	//   **  * 
        11'h6d7: data = 8'b00110010;	//   **  * 
        11'h6d8: data = 8'b00110010;	//   **  * 
        11'h6d9: data = 8'b00100010;	//   *   * 
        11'h6da: data = 8'b00000000;	//         
        11'h6db: data = 8'b00000000;	//         
        11'h6dc: data = 8'b00000000;	//         
        11'h6dd: data = 8'b00000000;	//         
        11'h6de: data = 8'b00000000;	//         
        11'h6df: data = 8'b00000000;	//         

    // code x6e (ื)
        11'he370: data = 8'b00000000;
        11'he371: data = 8'b00000000;
        11'he372: data = 8'b00010100;
        11'he373: data = 8'b00010100;
        11'he374: data = 8'b00111100;
        11'he375: data = 8'b01000010;
        11'he376: data = 8'b01111110;
        11'he377: data = 8'b00000000;
        11'he378: data = 8'b00000000;
        11'he379: data = 8'b00000000;
        11'he37a: data = 8'b00000000;
        11'he37b: data = 8'b00000000;
        11'he37c: data = 8'b00000000;
        11'he37d: data = 8'b00000000;
        11'he37e: data = 8'b00000000;
        11'he37f: data = 8'b00000000;

    // code x6f (น)
        11'h6f0: data = 8'b00000000;	//         
        11'h6f1: data = 8'b00000000;	//         
        11'h6f2: data = 8'b00000000;	//         
        11'h6f3: data = 8'b01100010;	//  **   * 
        11'h6f4: data = 8'b01100010;	//  **   * 
        11'h6f5: data = 8'b00100010;	//   *   * 
        11'h6f6: data = 8'b00100010;	//   *   * 
        11'h6f7: data = 8'b00100110;	//   *  ** 
        11'h6f8: data = 8'b00111010;	//   *** * 
        11'h6f9: data = 8'b00110110;	//   ** ** 
        11'h6fa: data = 8'b00000000;	//         
        11'h6fb: data = 8'b00000000;	//         
        11'h6fc: data = 8'b00000000;	//         
        11'h6fd: data = 8'b00000000;	//         
        11'h6fe: data = 8'b00000000;	//         
        11'h6ff: data = 8'b00000000;	//         

    // code x70 (ย)
        11'h700: data = 8'b00000000;	//         
        11'h701: data = 8'b00000000;	//         
        11'h702: data = 8'b00000000;	//         
        11'h703: data = 8'b01100100;	//  **  *  
        11'h704: data = 8'b01100100;	//  **  *  
        11'h705: data = 8'b01000100;	//  *   *  
        11'h706: data = 8'b01110100;	//  *** *  
        11'h707: data = 8'b01000100;	//  *   *  
        11'h708: data = 8'b01000100;	//  *   *  
        11'h709: data = 8'b00111000;	//   ***   
        11'h70a: data = 8'b00000000;	//         
        11'h70b: data = 8'b00000000;	//         
        11'h70c: data = 8'b00000000;	//         
        11'h70d: data = 8'b00000000;	//         
        11'h70e: data = 8'b00000000;	//         
        11'h70f: data = 8'b00000000;	//         

    // code x71 (ๆ)
        11'h710: data = 8'b00000000;	//         
        11'h711: data = 8'b00000000;	//         
        11'h712: data = 8'b00000000;	//         
        11'h713: data = 8'b00101000;	//   * *   
        11'h714: data = 8'b01010100;	//  * * *  
        11'h715: data = 8'b01100100;	//  **  *  
        11'h716: data = 8'b01110100;	//  *** *  
        11'h717: data = 8'b01100100;	//  **  *  
        11'h718: data = 8'b00000100;	//      *  
        11'h719: data = 8'b00000100;	//      *  
        11'h71a: data = 8'b00000100;	//      *  
        11'h71b: data = 8'b00000100;	//      *  
        11'h71c: data = 8'b00000100;	//      *  
        11'h71d: data = 8'b00000000;	//         
        11'h71e: data = 8'b00000000;	//         
        11'h71f: data = 8'b00000000;	//         

    // code x72 (พ)
        11'h720: data = 8'b00000000;	//         
        11'h721: data = 8'b00000000;	//         
        11'h722: data = 8'b00000000;	//         
        11'h723: data = 8'b01101101;	//  ** ** *
        11'h724: data = 8'b00101101;	//   * ** *
        11'h725: data = 8'b01101101;	//  ** ** *
        11'h726: data = 8'b00110011;	//   **  **
        11'h727: data = 8'b00110011;	//   **  **
        11'h728: data = 8'b00110011;	//   **  **
        11'h729: data = 8'b00100001;	//   *    *
        11'h72a: data = 8'b00000000;	//         
        11'h72b: data = 8'b00000000;	//         
        11'h72c: data = 8'b00000000;	//         
        11'h72d: data = 8'b00000000;	//         
        11'h72e: data = 8'b00000000;	//         
        11'h72f: data = 8'b00000000;	//         

    // code x73 (ห)
        11'h730: data = 8'b00000000;	//         
        11'h731: data = 8'b00000000;	//         
        11'h732: data = 8'b00000000;	//         
        11'h733: data = 8'b01100100;	//  **  *  
        11'h734: data = 8'b00100010;	//   *   * 
        11'h735: data = 8'b01100110;	//  **  ** 
        11'h736: data = 8'b00101010;	//   * * * 
        11'h737: data = 8'b00111010;	//   *** * 
        11'h738: data = 8'b00110010;	//   **  * 
        11'h739: data = 8'b00100010;	//   *   * 
        11'h73a: data = 8'b00000000;	//         
        11'h73b: data = 8'b00000000;	//         
        11'h73c: data = 8'b00000000;	//         
        11'h73d: data = 8'b00000000;	//         
        11'h73e: data = 8'b00000000;	//         
        11'h73f: data = 8'b00000000;	//         

    // code x74 (ะ)
        11'h740: data = 8'b00000000;	//         
        11'h741: data = 8'b00000000;	//         
        11'h742: data = 8'b00000000;	//         
        11'h743: data = 8'b01101000;	//  ** *   
        11'h744: data = 8'b11111000;	// *****   
        11'h745: data = 8'b01110000;	//  ***    
        11'h746: data = 8'b00000000;	//         
        11'h747: data = 8'b01101000;	//  ** *   
        11'h748: data = 8'b11111000;	// *****   
        11'h749: data = 8'b01110000;	//  ***    
        11'h74a: data = 8'b00000000;	//         
        11'h74b: data = 8'b00000000;	//         
        11'h74c: data = 8'b00000000;	//         
        11'h74d: data = 8'b00000000;	//         
        11'h74e: data = 8'b00000000;	//         
        11'h74f: data = 8'b00000000;	//         

    // code x75 (ี)
        11'he350: data = 8'b00000000;
        11'he351: data = 8'b00000000;
        11'he352: data = 8'b00000010;
        11'he353: data = 8'b00000010;
        11'he354: data = 8'b00111100;
        11'he355: data = 8'b01000010;
        11'he356: data = 8'b01111110;
        11'he357: data = 8'b00000000;
        11'he358: data = 8'b00000000;
        11'he359: data = 8'b00000000;
        11'he35a: data = 8'b00000000;
        11'he35b: data = 8'b00000000;
        11'he35c: data = 8'b00000000;
        11'he35d: data = 8'b00000000;
        11'he35e: data = 8'b00000000;
        11'he35f: data = 8'b00000000;

    // code x76 (อ)
        11'h760: data = 8'b00000000;	//         
        11'h761: data = 8'b00000000;	//         
        11'h762: data = 8'b00000000;	//         
        11'h763: data = 8'b01111000;	//  ****   
        11'h764: data = 8'b01000100;	//  *   *  
        11'h765: data = 8'b01100100;	//  **  *  
        11'h766: data = 8'b01010100;	//  * * *  
        11'h767: data = 8'b01100100;	//  **  *  
        11'h768: data = 8'b01000100;	//  *   *  
        11'h769: data = 8'b00111000;	//   ***   
        11'h76a: data = 8'b00000000;	//         
        11'h76b: data = 8'b00000000;	//         
        11'h76c: data = 8'b00000000;	//         
        11'h76d: data = 8'b00000000;	//         
        11'h76e: data = 8'b00000000;	//         
        11'h76f: data = 8'b00000000;	//         

    // code x77 (ไ)
        11'h770: data = 8'b10100000;	// * *     
        11'h771: data = 8'b00100000;	//   *     
        11'h772: data = 8'b00100000;	//   *     
        11'h773: data = 8'b00100000;	//   *     
        11'h774: data = 8'b00100000;	//   *     
        11'h775: data = 8'b00100000;	//   *     
        11'h776: data = 8'b00100000;	//   *     
        11'h777: data = 8'b00110000;	//   **    
        11'h778: data = 8'b00110000;	//   **    
        11'h779: data = 8'b00110000;	//   **    
        11'h77a: data = 8'b00000000;	//         
        11'h77b: data = 8'b00000000;	//         
        11'h77c: data = 8'b00000000;	//         
        11'h77d: data = 8'b00000000;	//         
        11'h77e: data = 8'b00000000;	//         
        11'h77f: data = 8'b00000000;	//         

    // code x78 (ป)
        11'h780: data = 8'b00000010;	//       * 
        11'h781: data = 8'b00000010;	//       * 
        11'h782: data = 8'b00000010;	//       * 
        11'h783: data = 8'b01100010;	//  **   * 
        11'h784: data = 8'b01100010;	//  **   * 
        11'h785: data = 8'b00100010;	//   *   * 
        11'h786: data = 8'b00100010;	//   *   * 
        11'h787: data = 8'b00100010;	//   *   * 
        11'h788: data = 8'b00100010;	//   *   * 
        11'h789: data = 8'b00011100;	//    ***  
        11'h78a: data = 8'b00000000;	//         
        11'h78b: data = 8'b00000000;	//         
        11'h78c: data = 8'b00000000;	//         
        11'h78d: data = 8'b00000000;	//         
        11'h78e: data = 8'b00000000;	//         
        11'h78f: data = 8'b00000000;	//         

    // code x79 (ั)
        11'h790: data = 8'b10000000;	// *       
        11'h791: data = 8'b00000000;	//         
        11'h792: data = 8'b00000000;	//         
        11'h793: data = 8'b00000000;	//         
        11'h794: data = 8'b00000000;	//         
        11'h795: data = 8'b00000000;	//         
        11'h796: data = 8'b00000000;	//         
        11'h797: data = 8'b00000000;	//         
        11'h798: data = 8'b00000000;	//         
        11'h799: data = 8'b00000000;	//         
        11'h79a: data = 8'b00000000;	//         
        11'h79b: data = 8'b00000000;	//         
        11'h79c: data = 8'b00000000;	//         
        11'h79d: data = 8'b00000000;	//         
        11'h79e: data = 8'b00000000;	//         
        11'h79f: data = 8'b00000000;	//         

    // code x7a (ผ)
        11'h7a0: data = 8'b00000000;	//         
        11'h7a1: data = 8'b00000000;	//         
        11'h7a2: data = 8'b00000000;	//         
        11'h7a3: data = 8'b01100100;	//  **  *  
        11'h7a4: data = 8'b01100100;	//  **  *  
        11'h7a5: data = 8'b01100100;	//  **  *  
        11'h7a6: data = 8'b01000100;	//  *   *  
        11'h7a7: data = 8'b01010100;	//  * * *  
        11'h7a8: data = 8'b01101100;	//  ** **  
        11'h7a9: data = 8'b01000100;	//  *   *  
        11'h7aa: data = 8'b00000000;	//         
        11'h7ab: data = 8'b00000000;	//         
        11'h7ac: data = 8'b00000000;	//         
        11'h7ad: data = 8'b00000000;	//         
        11'h7ae: data = 8'b00000000;	//         
        11'h7af: data = 8'b00000000;	//         

    // code x41 (ฤ)
        11'h410: data = 8'b00000000;	//         
        11'h411: data = 8'b00000000;	//         
        11'h412: data = 8'b00000000;	//         
        11'h413: data = 8'b00111000;	//   ***   
        11'h414: data = 8'b01000100;	//  *   *  
        11'h415: data = 8'b01100100;	//  **  *  
        11'h416: data = 8'b01000100;	//  *   *  
        11'h417: data = 8'b01000100;	//  *   *  
        11'h418: data = 8'b01100100;	//  **  *  
        11'h419: data = 8'b01100100;	//  **  *  
        11'h41a: data = 8'b00000100;	//      *  
        11'h41b: data = 8'b00000100;	//      *  
        11'h41c: data = 8'b00000100;	//      *  
        11'h41d: data = 8'b00000000;	//         
        11'h41e: data = 8'b00000000;	//         
        11'h41f: data = 8'b00000000;	//         

    // code x42 (ฺ)
        11'h420: data = 8'b11111111;	// ********
        11'h421: data = 8'b11111111;	// ********
        11'h422: data = 8'b11111111;	// ********
        11'h423: data = 8'b11111111;	// ********
        11'h424: data = 8'b11111111;	// ********
        11'h425: data = 8'b11111111;	// ********
        11'h426: data = 8'b11111111;	// ********
        11'h427: data = 8'b11111111;	// ********
        11'h428: data = 8'b11111111;	// ********
        11'h429: data = 8'b11111111;	// ********
        11'h42a: data = 8'b11111111;	// ********
        11'h42b: data = 8'b11111111;	// ********
        11'h42c: data = 8'b11111111;	// ********
        11'h42d: data = 8'b11111111;	// ********
        11'h42e: data = 8'b11111111;	// ********
        11'h42f: data = 8'b11111111;	// ********

    // code x43 (ฉ)
        11'h430: data = 8'b00000000;	//         
        11'h431: data = 8'b00000000;	//         
        11'h432: data = 8'b00000000;	//         
        11'h433: data = 8'b01110000;	//  ***    
        11'h434: data = 8'b10001000;	// *   *   
        11'h435: data = 8'b11001000;	// **  *   
        11'h436: data = 8'b10001000;	// *   *   
        11'h437: data = 8'b11001000;	// **  *   
        11'h438: data = 8'b01111000;	//  ****   
        11'h439: data = 8'b01011000;	//  * **   
        11'h43a: data = 8'b00000000;	//         
        11'h43b: data = 8'b00000000;	//         
        11'h43c: data = 8'b00000000;	//         
        11'h43d: data = 8'b00000000;	//         
        11'h43e: data = 8'b00000000;	//         
        11'h43f: data = 8'b00000000;	//         

    // code x44 (ฏ)
        11'h440: data = 8'b00000000;	//         
        11'h441: data = 8'b00000000;	//         
        11'h442: data = 8'b00000000;	//         
        11'h443: data = 8'b00111000;	//   ***   
        11'h444: data = 8'b01100100;	//  **  *  
        11'h445: data = 8'b00100100;	//   *  *  
        11'h446: data = 8'b00100100;	//   *  *  
        11'h447: data = 8'b01100100;	//  **  *  
        11'h448: data = 8'b11000100;	// **   *  
        11'h449: data = 8'b01100100;	//  **  *  
        11'h44a: data = 8'b00000100;	//      *  
        11'h44b: data = 8'b01110100;	//  *** *  
        11'h44c: data = 8'b01111100;	//  *****  
        11'h44d: data = 8'b00000100;	//      *  
        11'h44e: data = 8'b00000000;	//         
        11'h44f: data = 8'b00000000;	//         

    // code x45 (ฎ)
        11'h450: data = 8'b00000000;	//         
        11'h451: data = 8'b00000000;	//         
        11'h452: data = 8'b00000000;	//         
        11'h453: data = 8'b00111000;	//   ***   
        11'h454: data = 8'b01100100;	//  **  *  
        11'h455: data = 8'b00100100;	//   *  *  
        11'h456: data = 8'b00100100;	//   *  *  
        11'h457: data = 8'b01100100;	//  **  *  
        11'h458: data = 8'b11000100;	// **   *  
        11'h459: data = 8'b01100100;	//  **  *  
        11'h45a: data = 8'b00000100;	//      *  
        11'h45b: data = 8'b00110100;	//   ** *  
        11'h45c: data = 8'b01111100;	//  *****  
        11'h45d: data = 8'b00100100;	//   *  *  
        11'h45e: data = 8'b00000000;	//         
        11'h45f: data = 8'b00000000;	//         

    // code x46 (โ)
        11'h460: data = 8'b11000000;	// **      
        11'h461: data = 8'b00100000;	//   *     
        11'h462: data = 8'b00100000;	//   *     
        11'h463: data = 8'b00100000;	//   *     
        11'h464: data = 8'b00100000;	//   *     
        11'h465: data = 8'b00100000;	//   *     
        11'h466: data = 8'b00100000;	//   *     
        11'h467: data = 8'b00110000;	//   **    
        11'h468: data = 8'b00100000;	//   *     
        11'h469: data = 8'b00110000;	//   **    
        11'h46a: data = 8'b00000000;	//         
        11'h46b: data = 8'b00000000;	//         
        11'h46c: data = 8'b00000000;	//         
        11'h46d: data = 8'b00000000;	//         
        11'h46e: data = 8'b00000000;	//         
        11'h46f: data = 8'b00000000;	//         

    // code x47 (ฌ)
        11'h470: data = 8'b00000000;	//         
        11'h471: data = 8'b00000000;	//         
        11'h472: data = 8'b00000000;	//         
        11'h473: data = 8'b00111001;	//   ***  *
        11'h474: data = 8'b01000101;	//  *   * *
        11'h475: data = 8'b01100101;	//  **  * *
        11'h476: data = 8'b01000101;	//  *   * *
        11'h477: data = 8'b01101101;	//  ** ** *
        11'h478: data = 8'b00100111;	//   *  ***
        11'h479: data = 8'b01101101;	//  ** ** *
        11'h47a: data = 8'b00000000;	//         
        11'h47b: data = 8'b00000000;	//         
        11'h47c: data = 8'b00000000;	//         
        11'h47d: data = 8'b00000000;	//         
        11'h47e: data = 8'b00000000;	//         
        11'h47f: data = 8'b00000000;	//         

    // code x48 (็)
        11'he580: data = 8'b00000000;
        11'he581: data = 8'b00000000;
        11'he582: data = 8'b00000010;
        11'he583: data = 8'b00000010;
        11'he584: data = 8'b00000010;
        11'he585: data = 8'b00111100;
        11'he586: data = 8'b01100110;
        11'he587: data = 8'b01010010;
        11'he588: data = 8'b01110110;
        11'he589: data = 8'b01101100;
        11'he58a: data = 8'b00000000;
        11'he58b: data = 8'b00000000;
        11'he58c: data = 8'b00000000;
        11'he58d: data = 8'b00000000;
        11'he58e: data = 8'b00000000;
        11'he58f: data = 8'b00000000;

    // code x49 (ณ)
        11'h490: data = 8'b00000000;	//         
        11'h491: data = 8'b00000000;	//         
        11'h492: data = 8'b00000000;	//         
        11'h493: data = 8'b00111000;	//   ***   
        11'h494: data = 8'b01000100;	//  *   *  
        11'h495: data = 8'b01100100;	//  **  *  
        11'h496: data = 8'b01000100;	//  *   *  
        11'h497: data = 8'b01100101;	//  **  * *
        11'h498: data = 8'b01110110;	//  *** ** 
        11'h499: data = 8'b01100101;	//  **  * *
        11'h49a: data = 8'b00000000;	//         
        11'h49b: data = 8'b00000000;	//         
        11'h49c: data = 8'b00000000;	//         
        11'h49d: data = 8'b00000000;	//         
        11'h49e: data = 8'b00000000;	//         
        11'h49f: data = 8'b00000000;	//         

    // code x4a (๋)
        11'h4a0: data = 8'b00000000;
        11'h4a1: data = 8'b00000000;
        11'h4a2: data = 8'b00000000;
        11'h4a3: data = 8'b00000000;
        11'h4a4: data = 8'b00011000;
        11'h4a5: data = 8'b00011000;
        11'h4a6: data = 8'b01111110;
        11'h4a7: data = 8'b01111110;
        11'h4a8: data = 8'b00011000;
        11'h4a9: data = 8'b00011000;
        11'h4aa: data = 8'b00000000;
        11'h4ab: data = 8'b00000000;
        11'h4ac: data = 8'b00000000;
        11'h4ad: data = 8'b00000000;
        11'h4ae: data = 8'b00000000;
        11'h4af: data = 8'b00000000;

    // code x4b (ษ)
        11'h4b0: data = 8'b00000000;	//         
        11'h4b1: data = 8'b00000000;	//         
        11'h4b2: data = 8'b00000000;	//         
        11'h4b3: data = 8'b01100010;	//  **   * 
        11'h4b4: data = 8'b00100010;	//   *   * 
        11'h4b5: data = 8'b01101010;	//  ** * * 
        11'h4b6: data = 8'b00101110;	//   * *** 
        11'h4b7: data = 8'b00100010;	//   *   * 
        11'h4b8: data = 8'b00100010;	//   *   * 
        11'h4b9: data = 8'b00011100;	//    ***  
        11'h4ba: data = 8'b00000000;	//         
        11'h4bb: data = 8'b00000000;	//         
        11'h4bc: data = 8'b00000000;	//         
        11'h4bd: data = 8'b00000000;	//         
        11'h4be: data = 8'b00000000;	//         
        11'h4bf: data = 8'b00000000;	//         

    // code x4c (ศ)
        11'h4c0: data = 8'b00000000;	//         
        11'h4c1: data = 8'b00000000;	//         
        11'h4c2: data = 8'b00001000;	//     *   
        11'h4c3: data = 8'b01111000;	//  ****   
        11'h4c4: data = 8'b11011000;	// ** **   
        11'h4c5: data = 8'b10101000;	// * * *   
        11'h4c6: data = 8'b11101000;	// *** *   
        11'h4c7: data = 8'b11101000;	// *** *   
        11'h4c8: data = 8'b10001000;	// *   *   
        11'h4c9: data = 8'b10001000;	// *   *   
        11'h4ca: data = 8'b00000000;	//         
        11'h4cb: data = 8'b00000000;	//         
        11'h4cc: data = 8'b00000000;	//         
        11'h4cd: data = 8'b00000000;	//         
        11'h4ce: data = 8'b00000000;	//         
        11'h4cf: data = 8'b00000000;	//         

    // code x4d (?)
        11'h4d0: data = 8'b00000000;	//         
        11'h4d1: data = 8'b00000000;	//         
        11'h4d2: data = 8'b01110000;	//  ***    
        11'h4d3: data = 8'b00001000;	//     *   
        11'h4d4: data = 8'b00001000;	//     *   
        11'h4d5: data = 8'b00010000;	//    *    
        11'h4d6: data = 8'b00110000;	//   **    
        11'h4d7: data = 8'b00100000;	//   *     
        11'h4d8: data = 8'b00000000;	//         
        11'h4d9: data = 8'b00100000;	//   *     
        11'h4da: data = 8'b00000000;	//         
        11'h4db: data = 8'b00000000;	//         
        11'h4dc: data = 8'b00000000;	//         
        11'h4dd: data = 8'b00000000;	//         
        11'h4de: data = 8'b00000000;	//         
        11'h4df: data = 8'b00000000;	//         

    // code x4e (์)
        11'h4e0: data = 8'b00000000;	//         
        11'h4e1: data = 8'b00000000;	//         
        11'h4e2: data = 8'b00000000;	//         
        11'h4e3: data = 8'b00000000;	//         
        11'h4e4: data = 8'b00000000;	//         
        11'h4e5: data = 8'b00000000;	//         
        11'h4e6: data = 8'b00000000;	//         
        11'h4e7: data = 8'b00000000;	//         
        11'h4e8: data = 8'b00000000;	//         
        11'h4e9: data = 8'b00000000;	//         
        11'h4ea: data = 8'b00000000;	//         
        11'h4eb: data = 8'b00000000;	//         
        11'h4ec: data = 8'b00000000;	//         
        11'h4ed: data = 8'b00000000;	//         
        11'h4ee: data = 8'b00000000;	//         
        11'h4ef: data = 8'b00000000;	//         

    // code x4f (ฯ)
        11'h4f0: data = 8'b00000000;	//         
        11'h4f1: data = 8'b00000000;	//         
        11'h4f2: data = 8'b00000000;	//         
        11'h4f3: data = 8'b11011000;	// ** **   
        11'h4f4: data = 8'b10101000;	// * * *   
        11'h4f5: data = 8'b11101000;	// *** *   
        11'h4f6: data = 8'b00001000;	//     *   
        11'h4f7: data = 8'b00001000;	//     *   
        11'h4f8: data = 8'b00001000;	//     *   
        11'h4f9: data = 8'b00001000;	//     *   
        11'h4fa: data = 8'b00000000;	//         
        11'h4fb: data = 8'b00000000;	//         
        11'h4fc: data = 8'b00000000;	//         
        11'h4fd: data = 8'b00000000;	//         
        11'h4fe: data = 8'b00000000;	//         
        11'h4ff: data = 8'b00000000;	//         

    // code x50 (ญ)
        11'h500: data = 8'b00000000;	//         
        11'h501: data = 8'b00000000;	//         
        11'h502: data = 8'b00000000;	//         
        11'h503: data = 8'b01111000;	//  ****   
        11'h504: data = 8'b01000100;	//  *   *  
        11'h505: data = 8'b01100100;	//  **  *  
        11'h506: data = 8'b01000100;	//  *   *  
        11'h507: data = 8'b01100100;	//  **  *  
        11'h508: data = 8'b01110100;	//  *** *  
        11'h509: data = 8'b01100111;	//  **  ***
        11'h50a: data = 8'b00000110;	//      ** 
        11'h50b: data = 8'b00000110;	//      ** 
        11'h50c: data = 8'b00000011;	//       **
        11'h50d: data = 8'b00000000;	//         
        11'h50e: data = 8'b00000000;	//         
        11'h50f: data = 8'b00000000;	//         

    // code x51 (๐)
        11'h510: data = 8'b00000000;	//         
        11'h511: data = 8'b00000000;	//         
        11'h512: data = 8'b00000000;	//         
        11'h513: data = 8'b00000000;	//         
        11'h514: data = 8'b00000000;	//         
        11'h515: data = 8'b00111100;	//   ****  
        11'h516: data = 8'b01100110;	//  **  ** 
        11'h517: data = 8'b01000010;	//  *    * 
        11'h518: data = 8'b01100110;	//  **  ** 
        11'h519: data = 8'b00111100;	//   ****  
        11'h51a: data = 8'b00000000;	//         
        11'h51b: data = 8'b00000000;	//         
        11'h51c: data = 8'b00000000;	//         
        11'h51d: data = 8'b00000000;	//         
        11'h51e: data = 8'b00000000;	//         
        11'h51f: data = 8'b00000000;	//         

    // code x52 (ฑ)
        11'h520: data = 8'b00000000;	//         
        11'h521: data = 8'b00000000;	//         
        11'h522: data = 8'b00000000;	//         
        11'h523: data = 8'b01110110;	//  *** ** 
        11'h524: data = 8'b11011010;	// ** ** * 
        11'h525: data = 8'b10011010;	// *  ** * 
        11'h526: data = 8'b11111010;	// ***** * 
        11'h527: data = 8'b00110010;	//   **  * 
        11'h528: data = 8'b00110010;	//   **  * 
        11'h529: data = 8'b00100010;	//   *   * 
        11'h52a: data = 8'b00000000;	//         
        11'h52b: data = 8'b00000000;	//         
        11'h52c: data = 8'b00000000;	//         
        11'h52d: data = 8'b00000000;	//         
        11'h52e: data = 8'b00000000;	//         
        11'h52f: data = 8'b00000000;	//         

    // code x53 (ฆ)
        11'h530: data = 8'b00000000;	//         
        11'h531: data = 8'b00000000;	//         
        11'h532: data = 8'b00000000;	//         
        11'h533: data = 8'b01110100;	//  *** *  
        11'h534: data = 8'b11010100;	// ** * *  
        11'h535: data = 8'b10110100;	// * ** *  
        11'h536: data = 8'b11100100;	// ***  *  
        11'h537: data = 8'b01110100;	//  *** *  
        11'h538: data = 8'b01011100;	//  * ***  
        11'h539: data = 8'b01100100;	//  **  *  
        11'h53a: data = 8'b00000000;	//         
        11'h53b: data = 8'b00000000;	//         
        11'h53c: data = 8'b00000000;	//         
        11'h53d: data = 8'b00000000;	//         
        11'h53e: data = 8'b00000000;	//         
        11'h53f: data = 8'b00000000;	//         

    // code x54 (ธ)
        11'h540: data = 8'b00000000;	//         
        11'h541: data = 8'b00000000;	//         
        11'h542: data = 8'b00000000;	//         
        11'h543: data = 8'b01111000;	//  ****   
        11'h544: data = 8'b01100000;	//  **     
        11'h545: data = 8'b00011000;	//    **   
        11'h546: data = 8'b01001000;	//  *  *   
        11'h547: data = 8'b01001000;	//  *  *   
        11'h548: data = 8'b01001000;	//  *  *   
        11'h549: data = 8'b01111000;	//  ****   
        11'h54a: data = 8'b00000000;	//         
        11'h54b: data = 8'b00000000;	//         
        11'h54c: data = 8'b00000000;	//         
        11'h54d: data = 8'b00000000;	//         
        11'h54e: data = 8'b00000000;	//         
        11'h54f: data = 8'b00000000;	//         

    // code x55 (๊)
        11'he570: data = 8'b00000000;
        11'he571: data = 8'b00000000;
        11'he572: data = 8'b00000000;
        11'he573: data = 8'b00000001;
        11'he574: data = 8'b00000001;
        11'he575: data = 8'b00110111;
        11'he576: data = 8'b01001011;
        11'he577: data = 8'b01110011;
        11'he578: data = 8'b01110011;
        11'he579: data = 8'b00110010;
        11'he57a: data = 8'b00000000;
        11'he57b: data = 8'b00000000;
        11'he57c: data = 8'b00000000;
        11'he57d: data = 8'b00000000;
        11'he57e: data = 8'b00000000;
        11'he57f: data = 8'b00000000;

    // code x56 (ฮ)
        11'h560: data = 8'b00000000;	//         
        11'h561: data = 8'b00000000;	//         
        11'h562: data = 8'b00000000;	//         
        11'h563: data = 8'b01111100;	//  *****  
        11'h564: data = 8'b01111100;	//  *****  
        11'h565: data = 8'b01100100;	//  **  *  
        11'h566: data = 8'b01110100;	//  *** *  
        11'h567: data = 8'b01100100;	//  **  *  
        11'h568: data = 8'b01000100;	//  *   *  
        11'h569: data = 8'b00111000;	//   ***   
        11'h56a: data = 8'b00000000;	//         
        11'h56b: data = 8'b00000000;	//         
        11'h56c: data = 8'b00000000;	//         
        11'h56d: data = 8'b00000000;	//         
        11'h56e: data = 8'b00000000;	//         
        11'h56f: data = 8'b00000000;	//         

    // code x57 (")
        11'h570: data = 8'b00000000;	//         
        11'h571: data = 8'b00000000;	//         
        11'h572: data = 8'b01010000;	//  * *    
        11'h573: data = 8'b01010000;	//  * *    
        11'h574: data = 8'b01010000;	//  * *    
        11'h575: data = 8'b00000000;	//         
        11'h576: data = 8'b00000000;	//         
        11'h577: data = 8'b00000000;	//         
        11'h578: data = 8'b00000000;	//         
        11'h579: data = 8'b00000000;	//         
        11'h57a: data = 8'b00000000;	//         
        11'h57b: data = 8'b00000000;	//         
        11'h57c: data = 8'b00000000;	//         
        11'h57d: data = 8'b00000000;	//         
        11'h57e: data = 8'b00000000;	//         
        11'h57f: data = 8'b00000000;	//         

    // code x58 ())
        11'h580: data = 8'b00000000;	//         
        11'h581: data = 8'b00000000;	//         
        11'h582: data = 8'b01000000;	//  *      
        11'h583: data = 8'b01100000;	//  **     
        11'h584: data = 8'b00100000;	//   *     
        11'h585: data = 8'b00100000;	//   *     
        11'h586: data = 8'b00100000;	//   *     
        11'h587: data = 8'b00100000;	//   *     
        11'h588: data = 8'b00100000;	//   *     
        11'h589: data = 8'b01000000;	//  *      
        11'h58a: data = 8'b01000000;	//  *      
        11'h58b: data = 8'b00000000;	//         
        11'h58c: data = 8'b00000000;	//         
        11'h58d: data = 8'b00000000;	//         
        11'h58e: data = 8'b00000000;	//         
        11'h58f: data = 8'b00000000;	//         

    // code x59 (ํ)
        11'h590: data = 8'b11111111;	// ********
        11'h591: data = 8'b11111111;	// ********
        11'h592: data = 8'b11111111;	// ********
        11'h593: data = 8'b11111111;	// ********
        11'h594: data = 8'b11111111;	// ********
        11'h595: data = 8'b11111111;	// ********
        11'h596: data = 8'b11111111;	// ********
        11'h597: data = 8'b11111111;	// ********
        11'h598: data = 8'b11111111;	// ********
        11'h599: data = 8'b11111111;	// ********
        11'h59a: data = 8'b11111111;	// ********
        11'h59b: data = 8'b11111111;	// ********
        11'h59c: data = 8'b11111111;	// ********
        11'h59d: data = 8'b11111111;	// ********
        11'h59e: data = 8'b11111111;	// ********
        11'h59f: data = 8'b11111111;	// ********

    // code x5a (()
        11'h5a0: data = 8'b00000000;	//         
        11'h5a1: data = 8'b00000000;	//         
        11'h5a2: data = 8'b01000000;	//  *      
        11'h5a3: data = 8'b11000000;	// **      
        11'h5a4: data = 8'b10000000;	// *       
        11'h5a5: data = 8'b10000000;	// *       
        11'h5a6: data = 8'b10000000;	// *       
        11'h5a7: data = 8'b10000000;	// *       
        11'h5a8: data = 8'b10000000;	// *       
        11'h5a9: data = 8'b01000000;	//  *      
        11'h5aa: data = 8'b01000000;	//  *      
        11'h5ab: data = 8'b00000000;	//         
        11'h5ac: data = 8'b00000000;	//         
        11'h5ad: data = 8'b00000000;	//         
        11'h5ae: data = 8'b00000000;	//         
        11'h5af: data = 8'b00000000;	//         

    // code x30 (จ)
        11'h300: data = 8'b00000000;	//         
        11'h301: data = 8'b00000000;	//         
        11'h302: data = 8'b00000000;	//         
        11'h303: data = 8'b01110000;	//  ***    
        11'h304: data = 8'b10001000;	// *   *   
        11'h305: data = 8'b01001000;	//  *  *   
        11'h306: data = 8'b11101000;	// *** *   
        11'h307: data = 8'b01101000;	//  ** *   
        11'h308: data = 8'b00101000;	//   * *   
        11'h309: data = 8'b00111000;	//   ***   
        11'h30a: data = 8'b00000000;	//         
        11'h30b: data = 8'b00000000;	//         
        11'h30c: data = 8'b00000000;	//         
        11'h30d: data = 8'b00000000;	//         
        11'h30e: data = 8'b00000000;	//         
        11'h30f: data = 8'b00000000;	//         

    // code x31 (1)
        11'h310: data = 8'b00000000;	//         
        11'h311: data = 8'b00000000;	//         
        11'h312: data = 8'b00010000;	//    *    
        11'h313: data = 8'b00110000;	//   **    
        11'h314: data = 8'b00010000;	//    *    
        11'h315: data = 8'b00010000;	//    *    
        11'h316: data = 8'b00010000;	//    *    
        11'h317: data = 8'b00010000;	//    *    
        11'h318: data = 8'b00010000;	//    *    
        11'h319: data = 8'b00111000;	//   ***   
        11'h31a: data = 8'b00000000;	//         
        11'h31b: data = 8'b00000000;	//         
        11'h31c: data = 8'b00000000;	//         
        11'h31d: data = 8'b00000000;	//         
        11'h31e: data = 8'b00000000;	//         
        11'h31f: data = 8'b00000000;	//         

    // code x32 (/)
        11'h320: data = 8'b00000000;	//         
        11'h321: data = 8'b00000000;	//         
        11'h322: data = 8'b00001000;	//     *   
        11'h323: data = 8'b00010000;	//    *    
        11'h324: data = 8'b00010000;	//    *    
        11'h325: data = 8'b00100000;	//   *     
        11'h326: data = 8'b00100000;	//   *     
        11'h327: data = 8'b01000000;	//  *      
        11'h328: data = 8'b01000000;	//  *      
        11'h329: data = 8'b11000000;	// **      
        11'h32a: data = 8'b10000000;	// *       
        11'h32b: data = 8'b00000000;	//         
        11'h32c: data = 8'b00000000;	//         
        11'h32d: data = 8'b00000000;	//         
        11'h32e: data = 8'b00000000;	//         
        11'h32f: data = 8'b00000000;	//         

    // code x33 (-)
        11'h330: data = 8'b00000000;	//         
        11'h331: data = 8'b00000000;	//         
        11'h332: data = 8'b00000000;	//         
        11'h333: data = 8'b00000000;	//         
        11'h334: data = 8'b00000000;	//         
        11'h335: data = 8'b00000000;	//         
        11'h336: data = 8'b11100000;	// ***     
        11'h337: data = 8'b00000000;	//         
        11'h338: data = 8'b00000000;	//         
        11'h339: data = 8'b00000000;	//         
        11'h33a: data = 8'b00000000;	//         
        11'h33b: data = 8'b00000000;	//         
        11'h33c: data = 8'b00000000;	//         
        11'h33d: data = 8'b00000000;	//         
        11'h33e: data = 8'b00000000;	//         
        11'h33f: data = 8'b00000000;	//         

    // code x34 (ภ)
        11'h340: data = 8'b00000000;	//         
        11'h341: data = 8'b00000000;	//         
        11'h342: data = 8'b00000000;	//         
        11'h343: data = 8'b00111100;	//   ****  
        11'h344: data = 8'b00100010;	//   *   * 
        11'h345: data = 8'b01110010;	//  ***  * 
        11'h346: data = 8'b00100010;	//   *   * 
        11'h347: data = 8'b00100010;	//   *   * 
        11'h348: data = 8'b01100010;	//  **   * 
        11'h349: data = 8'b01100010;	//  **   * 
        11'h34a: data = 8'b00000000;	//         
        11'h34b: data = 8'b00000000;	//         
        11'h34c: data = 8'b00000000;	//         
        11'h34d: data = 8'b00000000;	//         
        11'h34e: data = 8'b00000000;	//         
        11'h34f: data = 8'b00000000;	//         

    // code x35 (ถ)
        11'h350: data = 8'b00000000;	//         
        11'h351: data = 8'b00000000;	//         
        11'h352: data = 8'b00000000;	//         
        11'h353: data = 8'b00111000;	//   ***   
        11'h354: data = 8'b01000100;	//  *   *  
        11'h355: data = 8'b01100100;	//  **  *  
        11'h356: data = 8'b01000100;	//  *   *  
        11'h357: data = 8'b01000100;	//  *   *  
        11'h358: data = 8'b01100100;	//  **  *  
        11'h359: data = 8'b01100100;	//  **  *  
        11'h35a: data = 8'b00000000;	//         
        11'h35b: data = 8'b00000000;	//         
        11'h35c: data = 8'b00000000;	//         
        11'h35d: data = 8'b00000000;	//         
        11'h35e: data = 8'b00000000;	//         
        11'h35f: data = 8'b00000000;	//         

    // code x36 (ุ)
        11'he380: data = 8'b00000000;
        11'he381: data = 8'b00000000;
        11'he382: data = 8'b00000000;
        11'he383: data = 8'b00000000;
        11'he384: data = 8'b00000000;
        11'he385: data = 8'b00000000;
        11'he386: data = 8'b00000000;
        11'he387: data = 8'b00000000;
        11'he388: data = 8'b00000000;
        11'he389: data = 8'b00010000;
        11'he38a: data = 8'b00101000;
        11'he38b: data = 8'b00011000;
        11'he38c: data = 8'b00001000;
        11'he38d: data = 8'b00001000;
        11'he38e: data = 8'b00000000;
        11'he38f: data = 8'b00000000;

    // code x37 (ึ)
        11'he360: data = 8'b00000000;
        11'he361: data = 8'b00000000;
        11'he362: data = 8'b00001100;
        11'he363: data = 8'b00001100;
        11'he364: data = 8'b00111110;
        11'he365: data = 8'b01000010;
        11'he366: data = 8'b01111110;
        11'he367: data = 8'b00000000;
        11'he368: data = 8'b00000000;
        11'he369: data = 8'b00000000;
        11'he36a: data = 8'b00000000;
        11'he36b: data = 8'b00000000;
        11'he36c: data = 8'b00000000;
        11'he36d: data = 8'b00000000;
        11'he36e: data = 8'b00000000;
        11'he36f: data = 8'b00000000;

    // code x38 (ค)
        11'h380: data = 8'b00000000;	//         
        11'h381: data = 8'b00000000;	//         
        11'h382: data = 8'b00000000;	//         
        11'h383: data = 8'b01110000;	//  ***    
        11'h384: data = 8'b11001000;	// **  *   
        11'h385: data = 8'b10101000;	// * * *   
        11'h386: data = 8'b11101000;	// *** *   
        11'h387: data = 8'b11101000;	// *** *   
        11'h388: data = 8'b10001000;	// *   *   
        11'h389: data = 8'b10001000;	// *   *   
        11'h38a: data = 8'b00000000;	//         
        11'h38b: data = 8'b00000000;	//         
        11'h38c: data = 8'b00000000;	//         
        11'h38d: data = 8'b00000000;	//         
        11'h38e: data = 8'b00000000;	//         
        11'h38f: data = 8'b00000000;	//         

    // code x39 (ต)
        11'h390: data = 8'b00000000;	//         
        11'h391: data = 8'b00000000;	//         
        11'h392: data = 8'b00000000;	//         
        11'h393: data = 8'b01111000;	//  ****   
        11'h394: data = 8'b10101000;	// * * *   
        11'h395: data = 8'b10101000;	// * * *   
        11'h396: data = 8'b10101000;	// * * *   
        11'h397: data = 8'b10101000;	// * * *   
        11'h398: data = 8'b11001000;	// **  *   
        11'h399: data = 8'b11001000;	// **  *   
        11'h39a: data = 8'b00000000;	//         
        11'h39b: data = 8'b00000000;	//         
        11'h39c: data = 8'b00000000;	//         
        11'h39d: data = 8'b00000000;	//         
        11'h39e: data = 8'b00000000;	//         
        11'h39f: data = 8'b00000000;	//         

    // code x21 (!)
        11'h210: data = 8'b00000000;	//         
        11'h211: data = 8'b00000000;	//         
        11'h212: data = 8'b01000000;	//  *      
        11'h213: data = 8'b01000000;	//  *      
        11'h214: data = 8'b01000000;	//  *      
        11'h215: data = 8'b01000000;	//  *      
        11'h216: data = 8'b01000000;	//  *      
        11'h217: data = 8'b01000000;	//  *      
        11'h218: data = 8'b01000000;	//  *      
        11'h219: data = 8'b01000000;	//  *      
        11'h21a: data = 8'b00000000;	//         
        11'h21b: data = 8'b00000000;	//         
        11'h21c: data = 8'b00000000;	//         
        11'h21d: data = 8'b00000000;	//         
        11'h21e: data = 8'b00000000;	//         
        11'h21f: data = 8'b00000000;	//         

    // code x22 (.)
        11'h220: data = 8'b00000000;	//         
        11'h221: data = 8'b00000000;	//         
        11'h222: data = 8'b00000000;	//         
        11'h223: data = 8'b00000000;	//         
        11'h224: data = 8'b00000000;	//         
        11'h225: data = 8'b00000000;	//         
        11'h226: data = 8'b00000000;	//         
        11'h227: data = 8'b00000000;	//         
        11'h228: data = 8'b01000000;	//  *      
        11'h229: data = 8'b01000000;	//  *      
        11'h22a: data = 8'b00000000;	//         
        11'h22b: data = 8'b00000000;	//         
        11'h22c: data = 8'b00000000;	//         
        11'h22d: data = 8'b00000000;	//         
        11'h22e: data = 8'b00000000;	//         
        11'h22f: data = 8'b00000000;	//         

    // code x23 (๒)
        11'h230: data = 8'b00000000;	//         
        11'h231: data = 8'b00000000;	//         
        11'h232: data = 8'b00000000;	//         
        11'h233: data = 8'b01000000;	//  *      
        11'h234: data = 8'b01000000;	//  *      
        11'h235: data = 8'b01011110;	//  * **** 
        11'h236: data = 8'b01111010;	//  **** * 
        11'h237: data = 8'b01010010;	//  * *  * 
        11'h238: data = 8'b01000010;	//  *    * 
        11'h239: data = 8'b00111100;	//   ****  
        11'h23a: data = 8'b00000000;	//         
        11'h23b: data = 8'b00000000;	//         
        11'h23c: data = 8'b00000000;	//         
        11'h23d: data = 8'b00000000;	//         
        11'h23e: data = 8'b00000000;	//         
        11'h23f: data = 8'b00000000;	//         

    // code x24 (๓)
        11'h240: data = 8'b00000000;	//         
        11'h241: data = 8'b00000000;	//         
        11'h242: data = 8'b00000000;	//         
        11'h243: data = 8'b00000000;	//         
        11'h244: data = 8'b00000000;	//         
        11'h245: data = 8'b00110110;	//   ** ** 
        11'h246: data = 8'b01001010;	//  *  * * 
        11'h247: data = 8'b01001010;	//  *  * * 
        11'h248: data = 8'b01101010;	//  ** * * 
        11'h249: data = 8'b00101010;	//   * * * 
        11'h24a: data = 8'b00000000;	//         
        11'h24b: data = 8'b00000000;	//         
        11'h24c: data = 8'b00000000;	//         
        11'h24d: data = 8'b00000000;	//         
        11'h24e: data = 8'b00000000;	//         
        11'h24f: data = 8'b00000000;	//         

    // code x25 (๔)
        11'h250: data = 8'b00000000;	//         
        11'h251: data = 8'b00000000;	//         
        11'h252: data = 8'b00000001;	//        *
        11'h253: data = 8'b00000001;	//        *
        11'h254: data = 8'b00000011;	//       **
        11'h255: data = 8'b00111110;	//   ***** 
        11'h256: data = 8'b01111000;	//  ****   
        11'h257: data = 8'b01011100;	//  * ***  
        11'h258: data = 8'b01001100;	//  *  **  
        11'h259: data = 8'b00111111;	//   ******
        11'h25a: data = 8'b00000000;	//         
        11'h25b: data = 8'b00000000;	//         
        11'h25c: data = 8'b00000000;	//         
        11'h25d: data = 8'b00000000;	//         
        11'h25e: data = 8'b00000000;	//         
        11'h25f: data = 8'b00000000;	//         

    // code x26 (฿)
        11'h260: data = 8'b00000000;	//         
        11'h261: data = 8'b00010000;	//    *    
        11'h262: data = 8'b01111000;	//  ****   
        11'h263: data = 8'b01000100;	//  *   *  
        11'h264: data = 8'b01000100;	//  *   *  
        11'h265: data = 8'b01111000;	//  ****   
        11'h266: data = 8'b01000100;	//  *   *  
        11'h267: data = 8'b01000100;	//  *   *  
        11'h268: data = 8'b01000100;	//  *   *  
        11'h269: data = 8'b01111000;	//  ****   
        11'h26a: data = 8'b00010000;	//    *    
        11'h26b: data = 8'b00000000;	//         
        11'h26c: data = 8'b00000000;	//         
        11'h26d: data = 8'b00000000;	//         
        11'h26e: data = 8'b00000000;	//         
        11'h26f: data = 8'b00000000;	//         

    // code x27 (ง)
        11'h270: data = 8'b00000000;	//         
        11'h271: data = 8'b00000000;	//         
        11'h272: data = 8'b00000000;	//         
        11'h273: data = 8'b00110000;	//   **    
        11'h274: data = 8'b01110000;	//  ***    
        11'h275: data = 8'b00110000;	//   **    
        11'h276: data = 8'b10010000;	// *  *    
        11'h277: data = 8'b11010000;	// ** *    
        11'h278: data = 8'b01110000;	//  ***    
        11'h279: data = 8'b00110000;	//   **    
        11'h27a: data = 8'b00000000;	//         
        11'h27b: data = 8'b00000000;	//         
        11'h27c: data = 8'b00000000;	//         
        11'h27d: data = 8'b00000000;	//         
        11'h27e: data = 8'b00000000;	//         
        11'h27f: data = 8'b00000000;	//         

    // code x28 (๖)
        11'h280: data = 8'b00000000;	//         
        11'h281: data = 8'b00000000;	//         
        11'h282: data = 8'b00000000;	//         
        11'h283: data = 8'b11000000;	// **      
        11'h284: data = 8'b01000000;	//  *      
        11'h285: data = 8'b01111100;	//  *****  
        11'h286: data = 8'b01100110;	//  **  ** 
        11'h287: data = 8'b01100010;	//  **   * 
        11'h288: data = 8'b01110110;	//  *** ** 
        11'h289: data = 8'b00111100;	//   ****  
        11'h28a: data = 8'b00000000;	//         
        11'h28b: data = 8'b00000000;	//         
        11'h28c: data = 8'b00000000;	//         
        11'h28d: data = 8'b00000000;	//         
        11'h28e: data = 8'b00000000;	//         
        11'h28f: data = 8'b00000000;	//         

    // code x29 (๗)
        11'h290: data = 8'b00000000;	//         
        11'h291: data = 8'b00000000;	//         
        11'h292: data = 8'b00000000;	//         
        11'h293: data = 8'b00000001;	//        *
        11'h294: data = 8'b00000001;	//        *
        11'h295: data = 8'b00110111;	//   ** ***
        11'h296: data = 8'b01001011;	//  *  * **
        11'h297: data = 8'b01110011;	//  ***  **
        11'h298: data = 8'b01110011;	//  ***  **
        11'h299: data = 8'b00110010;	//   **  * 
        11'h29a: data = 8'b00000000;	//         
        11'h29b: data = 8'b00000000;	//         
        11'h29c: data = 8'b00000000;	//         
        11'h29d: data = 8'b00000000;	//         
        11'h29e: data = 8'b00000000;	//         
        11'h29f: data = 8'b00000000;	//         

    // code x2a (๕)
        11'h2a0: data = 8'b00000000;	//         
        11'h2a1: data = 8'b00000000;	//         
        11'h2a2: data = 8'b00000001;	//        *
        11'h2a3: data = 8'b00011001;	//    **  *
        11'h2a4: data = 8'b00011110;	//    **** 
        11'h2a5: data = 8'b00111110;	//   ***** 
        11'h2a6: data = 8'b01110000;	//  ***    
        11'h2a7: data = 8'b01010000;	//  * *    
        11'h2a8: data = 8'b01011000;	//  * **   
        11'h2a9: data = 8'b00111110;	//   ***** 
        11'h2aa: data = 8'b00000000;	//         
        11'h2ab: data = 8'b00000000;	//         
        11'h2ac: data = 8'b00000000;	//         
        11'h2ad: data = 8'b00000000;	//         
        11'h2ae: data = 8'b00000000;	//         
        11'h2af: data = 8'b00000000;	//         

    // code x2b (๙)
        11'h2b0: data = 8'b00000000;	//         
        11'h2b1: data = 8'b00000000;	//         
        11'h2b2: data = 8'b00000001;	//        *
        11'h2b3: data = 8'b00000001;	//        *
        11'h2b4: data = 8'b00000001;	//        *
        11'h2b5: data = 8'b00111111;	//   ******
        11'h2b6: data = 8'b01001100;	//  *  **  
        11'h2b7: data = 8'b01010100;	//  * * *  
        11'h2b8: data = 8'b01111110;	//  ****** 
        11'h2b9: data = 8'b00110010;	//   **  * 
        11'h2ba: data = 8'b00000000;	//         
        11'h2bb: data = 8'b00000000;	//         
        11'h2bc: data = 8'b00000000;	//         
        11'h2bd: data = 8'b00000000;	//         
        11'h2be: data = 8'b00000000;	//         
        11'h2bf: data = 8'b00000000;	//         

    // code x2c (ม)
        11'h2c0: data = 8'b00000000;	//         
        11'h2c1: data = 8'b00000000;	//         
        11'h2c2: data = 8'b00000000;	//         
        11'h2c3: data = 8'b01100100;	//  **  *  
        11'h2c4: data = 8'b10100100;	// * *  *  
        11'h2c5: data = 8'b01100100;	//  **  *  
        11'h2c6: data = 8'b00100100;	//   *  *  
        11'h2c7: data = 8'b01110100;	//  *** *  
        11'h2c8: data = 8'b10111100;	// * ****  
        11'h2c9: data = 8'b01101100;	//  ** **  
        11'h2ca: data = 8'b00000000;	//         
        11'h2cb: data = 8'b00000000;	//         
        11'h2cc: data = 8'b00000000;	//         
        11'h2cd: data = 8'b00000000;	//         
        11'h2ce: data = 8'b00000000;	//         
        11'h2cf: data = 8'b00000000;	//         

    // code x2d (ข)
        11'h2d0: data = 8'b00000000;	//         
        11'h2d1: data = 8'b00000000;	//         
        11'h2d2: data = 8'b00000000;	//         
        11'h2d3: data = 8'b01110100;	//  *** *  
        11'h2d4: data = 8'b11010100;	// ** * *  
        11'h2d5: data = 8'b11010100;	// ** * *  
        11'h2d6: data = 8'b00100100;	//   *  *  
        11'h2d7: data = 8'b00100100;	//   *  *  
        11'h2d8: data = 8'b00100100;	//   *  *  
        11'h2d9: data = 8'b00111100;	//   ****  
        11'h2da: data = 8'b00000000;	//         
        11'h2db: data = 8'b00000000;	//         
        11'h2dc: data = 8'b00000000;	//         
        11'h2dd: data = 8'b00000000;	//         
        11'h2de: data = 8'b00000000;	//         
        11'h2df: data = 8'b00000000;	//         

    // code x2e (ใ)
        11'h2e0: data = 8'b11000000;	// **      
        11'h2e1: data = 8'b11000000;	// **      
        11'h2e2: data = 8'b01000000;	//  *      
        11'h2e3: data = 8'b01000000;	//  *      
        11'h2e4: data = 8'b01000000;	//  *      
        11'h2e5: data = 8'b01000000;	//  *      
        11'h2e6: data = 8'b01000000;	//  *      
        11'h2e7: data = 8'b01100000;	//  **     
        11'h2e8: data = 8'b00110000;	//   **    
        11'h2e9: data = 8'b01100000;	//  **     
        11'h2ea: data = 8'b00000000;	//         
        11'h2eb: data = 8'b00000000;	//         
        11'h2ec: data = 8'b00000000;	//         
        11'h2ed: data = 8'b00000000;	//         
        11'h2ee: data = 8'b00000000;	//         
        11'h2ef: data = 8'b00000000;	//         

    // code x2f (ฝ)
        11'h2f0: data = 8'b00000100;	//      *  
        11'h2f1: data = 8'b00000100;	//      *  
        11'h2f2: data = 8'b00000100;	//      *  
        11'h2f3: data = 8'b01100100;	//  **  *  
        11'h2f4: data = 8'b01100100;	//  **  *  
        11'h2f5: data = 8'b01100100;	//  **  *  
        11'h2f6: data = 8'b01000100;	//  *   *  
        11'h2f7: data = 8'b01010100;	//  * * *  
        11'h2f8: data = 8'b01101100;	//  ** **  
        11'h2f9: data = 8'b01000100;	//  *   *  
        11'h2fa: data = 8'b00000000;	//         
        11'h2fb: data = 8'b00000000;	//         
        11'h2fc: data = 8'b00000000;	//         
        11'h2fd: data = 8'b00000000;	//         
        11'h2fe: data = 8'b00000000;	//         
        11'h2ff: data = 8'b00000000;	//         

    // code x3a (ซ)
        11'h3a0: data = 8'b00000000;	//         
        11'h3a1: data = 8'b00000000;	//         
        11'h3a2: data = 8'b00000100;	//      *  
        11'h3a3: data = 8'b11110100;	// **** *  
        11'h3a4: data = 8'b11011100;	// ** ***  
        11'h3a5: data = 8'b10110100;	// * ** *  
        11'h3a6: data = 8'b11100100;	// ***  *  
        11'h3a7: data = 8'b00100100;	//   *  *  
        11'h3a8: data = 8'b00100100;	//   *  *  
        11'h3a9: data = 8'b00111100;	//   ****  
        11'h3aa: data = 8'b00000000;	//         
        11'h3ab: data = 8'b00000000;	//         
        11'h3ac: data = 8'b00000000;	//         
        11'h3ad: data = 8'b00000000;	//         
        11'h3ae: data = 8'b00000000;	//         
        11'h3af: data = 8'b00000000;	//         

    // code x3b (ว)
        11'h3b0: data = 8'b00000000;	//         
        11'h3b1: data = 8'b00000000;	//         
        11'h3b2: data = 8'b00000000;	//         
        11'h3b3: data = 8'b01110000;	//  ***    
        11'h3b4: data = 8'b11001000;	// **  *   
        11'h3b5: data = 8'b00001000;	//     *   
        11'h3b6: data = 8'b00001000;	//     *   
        11'h3b7: data = 8'b00011000;	//    **   
        11'h3b8: data = 8'b00101000;	//   * *   
        11'h3b9: data = 8'b00011000;	//    **   
        11'h3ba: data = 8'b00000000;	//         
        11'h3bb: data = 8'b00000000;	//         
        11'h3bc: data = 8'b00000000;	//         
        11'h3bd: data = 8'b00000000;	//         
        11'h3be: data = 8'b00000000;	//         
        11'h3bf: data = 8'b00000000;	//         

    // code x3c (ฒ)
        11'h3c0: data = 8'b00000000;	//         
        11'h3c1: data = 8'b00000000;	//         
        11'h3c2: data = 8'b00000000;	//         
        11'h3c3: data = 8'b01110001;	//  ***   *
        11'h3c4: data = 8'b10001001;	// *   *  *
        11'h3c5: data = 8'b10101001;	// * * *  *
        11'h3c6: data = 8'b10101001;	// * * *  *
        11'h3c7: data = 8'b10101001;	// * * *  *
        11'h3c8: data = 8'b11011111;	// ** *****
        11'h3c9: data = 8'b11011001;	// ** **  *
        11'h3ca: data = 8'b00000000;	//         
        11'h3cb: data = 8'b00000000;	//         
        11'h3cc: data = 8'b00000000;	//         
        11'h3cd: data = 8'b00000000;	//         
        11'h3ce: data = 8'b00000000;	//         
        11'h3cf: data = 8'b00000000;	//         

    // code x3d (ช)
        11'h3d0: data = 8'b00000000;	//         
        11'h3d1: data = 8'b00000000;	//         
        11'h3d2: data = 8'b00000000;	//         
        11'h3d3: data = 8'b01110100;	//  *** *  
        11'h3d4: data = 8'b11011100;	// ** ***  
        11'h3d5: data = 8'b11010100;	// ** * *  
        11'h3d6: data = 8'b00100100;	//   *  *  
        11'h3d7: data = 8'b00100100;	//   *  *  
        11'h3d8: data = 8'b00100100;	//   *  *  
        11'h3d9: data = 8'b00111100;	//   ****  
        11'h3da: data = 8'b00000000;	//         
        11'h3db: data = 8'b00000000;	//         
        11'h3dc: data = 8'b00000000;	//         
        11'h3dd: data = 8'b00000000;	//         
        11'h3de: data = 8'b00000000;	//         
        11'h3df: data = 8'b00000000;	//         

    // code x3e (ฬ)
        11'h3e0: data = 8'b00000000;	//         
        11'h3e1: data = 8'b00000000;	//         
        11'h3e2: data = 8'b00000000;	//         
        11'h3e3: data = 8'b01100011;	//  **   **
        11'h3e4: data = 8'b00100011;	//   *   **
        11'h3e5: data = 8'b01100001;	//  **    *
        11'h3e6: data = 8'b00101101;	//   * ** *
        11'h3e7: data = 8'b00101101;	//   * ** *
        11'h3e8: data = 8'b00110011;	//   **  **
        11'h3e9: data = 8'b00100001;	//   *    *
        11'h3ea: data = 8'b00000000;	//         
        11'h3eb: data = 8'b00000000;	//         
        11'h3ec: data = 8'b00000000;	//         
        11'h3ed: data = 8'b00000000;	//         
        11'h3ee: data = 8'b00000000;	//         
        11'h3ef: data = 8'b00000000;	//         

    // code x3f (ฦ)
        11'h3f0: data = 8'b00000000;	//         
        11'h3f1: data = 8'b00000000;	//         
        11'h3f2: data = 8'b00000000;	//         
        11'h3f3: data = 8'b00111000;	//   ***   
        11'h3f4: data = 8'b00100100;	//   *  *  
        11'h3f5: data = 8'b00100100;	//   *  *  
        11'h3f6: data = 8'b00100100;	//   *  *  
        11'h3f7: data = 8'b00100100;	//   *  *  
        11'h3f8: data = 8'b01100100;	//  **  *  
        11'h3f9: data = 8'b01100100;	//  **  *  
        11'h3fa: data = 8'b00000100;	//      *  
        11'h3fb: data = 8'b00000100;	//      *  
        11'h3fc: data = 8'b00000100;	//      *  
        11'h3fd: data = 8'b00000000;	//         
        11'h3fe: data = 8'b00000000;	//         
        11'h3ff: data = 8'b00000000;	//         

    // code x40 (๑)
        11'h400: data = 8'b00000000;	//         
        11'h401: data = 8'b00000000;	//         
        11'h402: data = 8'b00000000;	//         
        11'h403: data = 8'b00000000;	//         
        11'h404: data = 8'b00111100;	//   ****  
        11'h405: data = 8'b01100110;	//  **  ** 
        11'h406: data = 8'b01011010;	//  * ** * 
        11'h407: data = 8'b01001010;	//  *  * * 
        11'h408: data = 8'b01011010;	//  * ** * 
        11'h409: data = 8'b00110110;	//   ** ** 
        11'h40a: data = 8'b00000000;	//         
        11'h40b: data = 8'b00000000;	//         
        11'h40c: data = 8'b00000000;	//         
        11'h40d: data = 8'b00000000;	//         
        11'h40e: data = 8'b00000000;	//         
        11'h40f: data = 8'b00000000;	//         

    // code x5b (บ)
        11'h5b0: data = 8'b00000000;	//         
        11'h5b1: data = 8'b00000000;	//         
        11'h5b2: data = 8'b00000000;	//         
        11'h5b3: data = 8'b01100010;	//  **   * 
        11'h5b4: data = 8'b01100010;	//  **   * 
        11'h5b5: data = 8'b00100010;	//   *   * 
        11'h5b6: data = 8'b00100010;	//   *   * 
        11'h5b7: data = 8'b00100010;	//   *   * 
        11'h5b8: data = 8'b00100010;	//   *   * 
        11'h5b9: data = 8'b00011100;	//    ***  
        11'h5ba: data = 8'b00000000;	//         
        11'h5bb: data = 8'b00000000;	//         
        11'h5bc: data = 8'b00000000;	//         
        11'h5bd: data = 8'b00000000;	//         
        11'h5be: data = 8'b00000000;	//         
        11'h5bf: data = 8'b00000000;	//         

    // code x5c (ฃ)
        11'h5c0: data = 8'b00000000;	//         
        11'h5c1: data = 8'b00000000;	//         
        11'h5c2: data = 8'b00000000;	//         
        11'h5c3: data = 8'b01110100;	//  *** *  
        11'h5c4: data = 8'b11010100;	// ** * *  
        11'h5c5: data = 8'b10010100;	// *  * *  
        11'h5c6: data = 8'b11100100;	// ***  *  
        11'h5c7: data = 8'b00100100;	//   *  *  
        11'h5c8: data = 8'b00100100;	//   *  *  
        11'h5c9: data = 8'b00111100;	//   ****  
        11'h5ca: data = 8'b00000000;	//         
        11'h5cb: data = 8'b00000000;	//         
        11'h5cc: data = 8'b00000000;	//         
        11'h5cd: data = 8'b00000000;	//         
        11'h5ce: data = 8'b00000000;	//         
        11'h5cf: data = 8'b00000000;	//         

    // code x5d (ล)
        11'h5d0: data = 8'b00000000;	//         
        11'h5d1: data = 8'b00000000;	//         
        11'h5d2: data = 8'b00000000;	//         
        11'h5d3: data = 8'b01111000;	//  ****   
        11'h5d4: data = 8'b01000100;	//  *   *  
        11'h5d5: data = 8'b00111100;	//   ****  
        11'h5d6: data = 8'b01000100;	//  *   *  
        11'h5d7: data = 8'b01000100;	//  *   *  
        11'h5d8: data = 8'b01100100;	//  **  *  
        11'h5d9: data = 8'b01100100;	//  **  *  
        11'h5da: data = 8'b00000000;	//         
        11'h5db: data = 8'b00000000;	//         
        11'h5dc: data = 8'b00000000;	//         
        11'h5dd: data = 8'b00000000;	//         
        11'h5de: data = 8'b00000000;	//         
        11'h5df: data = 8'b00000000;	//         

    // code x5e (ู)
        11'he390: data = 8'b00000000;
        11'he391: data = 8'b00000000;
        11'he392: data = 8'b00000000;
        11'he393: data = 8'b00000000;
        11'he394: data = 8'b00000000;
        11'he395: data = 8'b00000000;
        11'he396: data = 8'b00000000;
        11'he397: data = 8'b00000000;
        11'he398: data = 8'b00000000;
        11'he399: data = 8'b00010010;
        11'he39a: data = 8'b00101010;
        11'he39b: data = 8'b00011010;
        11'he39c: data = 8'b00001010;
        11'he39d: data = 8'b00001010;
        11'he39e: data = 8'b00000100;
        11'he39f: data = 8'b00000000;

    // code x5f (๘)
        11'h5f0: data = 8'b00000000;	//         
        11'h5f1: data = 8'b00000000;	//         
        11'h5f2: data = 8'b00000010;	//       * 
        11'h5f3: data = 8'b00000010;	//       * 
        11'h5f4: data = 8'b00000010;	//       * 
        11'h5f5: data = 8'b00111100;	//   ****  
        11'h5f6: data = 8'b01100110;	//  **  ** 
        11'h5f7: data = 8'b01010010;	//  * *  * 
        11'h5f8: data = 8'b01110110;	//  *** ** 
        11'h5f9: data = 8'b01101100;	//  ** **  
        11'h5fa: data = 8'b00000000;	//         
        11'h5fb: data = 8'b00000000;	//         
        11'h5fc: data = 8'b00000000;	//         
        11'h5fd: data = 8'b00000000;	//         
        11'h5fe: data = 8'b00000000;	//         
        11'h5ff: data = 8'b00000000;	//         

    // code x60 (_)
        11'h600: data = 8'b00000000;	//         
        11'h601: data = 8'b00000000;	//         
        11'h602: data = 8'b00000000;	//         
        11'h603: data = 8'b00000000;	//         
        11'h604: data = 8'b00000000;	//         
        11'h605: data = 8'b00000000;	//         
        11'h606: data = 8'b00000000;	//         
        11'h607: data = 8'b00000000;	//         
        11'h608: data = 8'b00000000;	//         
        11'h609: data = 8'b00000000;	//         
        11'h60a: data = 8'b00000000;	//         
        11'h60b: data = 8'b00000000;	//         
        11'h60c: data = 8'b00000000;	//         
        11'h60d: data = 8'b11110000;	// ****    
        11'h60e: data = 8'b00000000;	//         
        11'h60f: data = 8'b00000000;	//         

    // code x7b (ฐ)
        11'h7b0: data = 8'b00000000;	//         
        11'h7b1: data = 8'b00000000;	//         
        11'h7b2: data = 8'b00000000;	//         
        11'h7b3: data = 8'b01111000;	//  ****   
        11'h7b4: data = 8'b01110000;	//  ***    
        11'h7b5: data = 8'b01101000;	//  ** *   
        11'h7b6: data = 8'b00101000;	//   * *   
        11'h7b7: data = 8'b01101000;	//  ** *   
        11'h7b8: data = 8'b00101000;	//   * *   
        11'h7b9: data = 8'b00111000;	//   ***   
        11'h7ba: data = 8'b00101000;	//   * *   
        11'h7bb: data = 8'b00101000;	//   * *   
        11'h7bc: data = 8'b11111000;	// *****   
        11'h7bd: data = 8'b01001000;	//  *  *   
        11'h7be: data = 8'b00000000;	//         
        11'h7bf: data = 8'b00000000;	//         

    // code x7c (ฅ)
        11'h7c0: data = 8'b00000000;	//         
        11'h7c1: data = 8'b00000000;	//         
        11'h7c2: data = 8'b00000000;	//         
        11'h7c3: data = 8'b11111000;	// *****   
        11'h7c4: data = 8'b10001000;	// *   *   
        11'h7c5: data = 8'b10101000;	// * * *   
        11'h7c6: data = 8'b11101000;	// *** *   
        11'h7c7: data = 8'b11101000;	// *** *   
        11'h7c8: data = 8'b10001000;	// *   *   
        11'h7c9: data = 8'b10001000;	// *   *   
        11'h7ca: data = 8'b00000000;	//         
        11'h7cb: data = 8'b00000000;	//         
        11'h7cc: data = 8'b00000000;	//         
        11'h7cd: data = 8'b00000000;	//         
        11'h7ce: data = 8'b00000000;	//         
        11'h7cf: data = 8'b00000000;	//         

    // code x7d (,)
        11'h7d0: data = 8'b00000000;	//         
        11'h7d1: data = 8'b00000000;	//         
        11'h7d2: data = 8'b00000000;	//         
        11'h7d3: data = 8'b00000000;	//         
        11'h7d4: data = 8'b00000000;	//         
        11'h7d5: data = 8'b00000000;	//         
        11'h7d6: data = 8'b00000000;	//         
        11'h7d7: data = 8'b00000000;	//         
        11'h7d8: data = 8'b01000000;	//  *      
        11'h7d9: data = 8'b01000000;	//  *      
        11'h7da: data = 8'b01000000;	//  *      
        11'h7db: data = 8'b01000000;	//  *      
        11'h7dc: data = 8'b00000000;	//         
        11'h7dd: data = 8'b00000000;	//         
        11'h7de: data = 8'b00000000;	//         
        11'h7df: data = 8'b00000000;	//         

    // code x7e (%)
        11'h7e0: data = 8'b00000000;	//         
        11'h7e1: data = 8'b00000000;	//         
        11'h7e2: data = 8'b01100010;	//  **   * 
        11'h7e3: data = 8'b10010100;	// *  * *  
        11'h7e4: data = 8'b10010100;	// *  * *  
        11'h7e5: data = 8'b01101111;	//  ** ****
        11'h7e6: data = 8'b00001100;	//     **  
        11'h7e7: data = 8'b00010100;	//    * *  
        11'h7e8: data = 8'b00110100;	//   ** *  
        11'h7e9: data = 8'b00100011;	//   *   **
        11'h7ea: data = 8'b00000000;	//         
        11'h7eb: data = 8'b00000000;	//         
        11'h7ec: data = 8'b00000000;	//         
        11'h7ed: data = 8'b00000000;	//         
        11'h7ee: data = 8'b00000000;	//         
        11'h7ef: data = 8'b00000000;	//         

    // code x20 ( )
        11'h200: data = 8'b11111111;	// ********
        11'h201: data = 8'b11111111;	// ********
        11'h202: data = 8'b11111111;	// ********
        11'h203: data = 8'b11111111;	// ********
        11'h204: data = 8'b11111111;	// ********
        11'h205: data = 8'b11111111;	// ********
        11'h206: data = 8'b11111111;	// ********
        11'h207: data = 8'b11111111;	// ********
        11'h208: data = 8'b11111111;	// ********
        11'h209: data = 8'b11111111;	// ********
        11'h20a: data = 8'b11111111;	// ********
        11'h20b: data = 8'b11111111;	// ********
        11'h20c: data = 8'b11111111;	// ********
        11'h20d: data = 8'b11111111;	// ********
        11'h20e: data = 8'b11111111;	// ********
        11'h20f: data = 8'b11111111;	// ********

            default: data = 8'b00000000; // Default to zero
        endcase
    endmodule
    
